* D:\University of Hail\2019-2020\Second\EE203 Electronic\Lab\ElectronicExp\app file\Experiment-5\Experiment-5.sch

* Schematics Version 9.1 - Web Update 1
* Sun Mar 22 19:56:33 2020



** Analysis setup **
.tran 20ns 3ms
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Experiment-5.net"
.INC "Experiment-5.als"


.probe


.END
