* D:\University of Hail\2019-2020\Second\EE203 Electronic\Lab\ElectronicExp\app file\Experiment-5\Schematic5.1o.sch

* Schematics Version 9.1 - Web Update 1
* Sat Mar 21 15:01:28 2020



** Analysis setup **
.tran 20ns 3ms
.OP 
.STMLIB "Schematic5.1o.stl"


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic5.1o.net"
.INC "Schematic5.1o.als"


.probe


.END
